`timescale 1ns / 1ps

module ledControl(
    input clk, rst
    );
endmodule
